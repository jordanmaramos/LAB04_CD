library verilog;
use verilog.vl_types.all;
entity LAB04_vlg_vec_tst is
end LAB04_vlg_vec_tst;
