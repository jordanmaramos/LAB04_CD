library verilog;
use verilog.vl_types.all;
entity DECODER_LOGICO_vlg_vec_tst is
end DECODER_LOGICO_vlg_vec_tst;
